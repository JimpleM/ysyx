`include"ysyx_23060077_riscv_define.v"
module ysyx_23060077_riscv_lsu(
    input 	                            clk,
    input 	                            rst_n,    

    input  	    [`DATA_WIDTH-1:0]       src1,
    input  	    [`DATA_WIDTH-1:0]       src2,
    input       [`DATA_WIDTH-1:0]       imm,

    input       [`LSU_OPT_WIDTH-1:0]    lsu_opt,
    input       [2:0]                   funct3,

    output                              mem_stall,
    output                              lsu_rd_wen,
    output  	  [`DATA_WIDTH-1:0]       lsu_result
);
wire ren;
wire wen;
wire [`DATA_WIDTH-1:0] raddr;
wire [`DATA_WIDTH-1:0] rdata;
wire [`DATA_WIDTH-1:0] waddr;
wire [`DATA_WIDTH-1:0] wdata;
wire [`DATA_WIDTH-1:0] wmask;
wire [`DATA_WIDTH-1:0]  mask;

wire [`DATA_WIDTH-1:0] rdata_t;
reg  [`DATA_WIDTH-1:0] rdata_r;
assign rdata = rdata_r;

reg wen_t;

assign mem_stall = ren | wen;

assign ren = (lsu_opt == `LSU_OPT_LOAD);
assign wen = (lsu_opt == `LSU_OPT_STORE);
assign raddr = src1 + imm;
assign waddr = src1 + imm;
assign wdata = src2;
assign wmask = mask;

ysyx_23060077_riscv_mux#(
    .NR_KEY      (5), 
    .KEY_LEN     (`LSU_OPT_WIDTH+3), 
    .DATA_LEN    (`DATA_WIDTH)
)riscv_mux_ls_lsu_opt(
  .key              ({lsu_opt,funct3}),
  .default_out      (0),
  .out              ({lsu_result}),
  .lut({{`LSU_OPT_LOAD,3'b000}, {{(`DATA_WIDTH-8){rdata[7]}}    ,rdata[7:0]},       //lb
        {`LSU_OPT_LOAD,3'b001}, {{(`DATA_WIDTH-16){rdata[15]}}  ,rdata[15:0]},      //lh
        {`LSU_OPT_LOAD,3'b010}, {{(`DATA_WIDTH-32){rdata[31]}}  ,rdata[31:0]},      //lw
        {`LSU_OPT_LOAD,3'b100}, {{(`DATA_WIDTH-8){1'b0}}        ,rdata[7:0]},       //lbu
        {`LSU_OPT_LOAD,3'b101}, {{(`DATA_WIDTH-16){1'b0}}       ,rdata[15:0]}       //lhu
  })
);


ysyx_23060077_riscv_mux#(
    .NR_KEY      (3), 
    .KEY_LEN     (`LSU_OPT_WIDTH+3), 
    .DATA_LEN    (`DATA_WIDTH)
)riscv_mux_ls_wmask(
  .key              ({lsu_opt,funct3}),
  .default_out      (0),
  .out              ({mask}),
  .lut({{`LSU_OPT_STORE,3'b000}, {32'd1},         //sb
        {`LSU_OPT_STORE,3'b001}, {32'd2},         //sh
        {`LSU_OPT_STORE,3'b010}, {32'd4}          //sw
  })
);


always @(posedge clk ) begin
  if(!rst_n)begin
    rdata_r <= 'd0;
  end
  else if(ren) begin
    rdata_r <= rdata_t;
  end
  else begin
    rdata_r <= 'd0;
  end
end

always @(posedge clk ) begin
  if(!rst_n)begin
    wen_t <= 'd0;
  end
  else if(wen) begin
    wen_t <= 'd1;
  end
  else begin
    wen_t <= 'd0;
  end
end
assign lsu_rd_wen = ren | wen;

// sim
import "DPI-C" function void riscv_pmem_read(input int raddr, output int rdata, input ren);
import "DPI-C" function void riscv_pmem_write(input int waddr, input int wdata,  input int wmask, input wen);

always @(*)begin
    riscv_pmem_read(raddr,rdata_t,ren);
    riscv_pmem_write(waddr,wdata,wmask,wen_t);
end

// ysyx_23060077_riscv_axi_lite  u_ysyx_23060077_riscv_axi_lite (
//     .aclk                   ( clk                                  ),
//     .areset_n               ( rst_n                                ),

//     .cpu_r_valid_i          (cpu_r_valid_i),
//     .cpu_r_addr_i           (raddr),
//     .cpu_r_ready_o          (cpu_r_ready_o),
//     .cpu_r_data_o           (inst),

//     .cpu_w_valid_i          (),
//     .cpu_w_addr_i           (),
//     .cpu_w_ready_o          (),
//     .cpu_w_data_i           (),
//     .cpu_w_strb_i           ()
// );


endmodule
