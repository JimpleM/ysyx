`include"ysyx_23060077_define.v"
`include"ysyx_23060077_axi_define.v"

module ysyx_23060077_Icache(
    input                       clock               ,
	input                       reset               ,
);

localparam b = 4;
localparam k = 16;




endmodule