
module ysyx_23060077_booth_code(
  
);


endmodule
