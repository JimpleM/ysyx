module riscv_sys_inst #(
    INST_WIDTH = 32,
    DATA_WIDTH = 32
) (
    input 	    [INPUT_WIDTH-1:0]       inst,
    output reg 	                        interrupt_status
);



endmodule